module (fie)
endmodule
